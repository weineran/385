module data_path
(
    input logic Clk, Reset, ClearA_LoadB, Run,
    input logic [7:0] switches,

)




