module adder2
(	
	input [1:0] A, B, 
	input Cin,
	output [1:0] S,
	output Cout
);

// Internal carries in the 2-bit adder				
wire c1;
full_adder FA0
(
	.x(A[0]), 
	.y(B[0]), 
	.z(Cin), 
	.s(S[0]), 
	.c(c1)
);
full_adder FA1
(
	.x(A[1]), 
	.y(B[1]), 
	.z(c1),  
	.s(S[1]), 
	.c(Cout)
);
	
endmodule
